
`ifndef ALU_VH
`define ALU_VH


`define ALU_NOP    5'b00000
`define ALU_SUM_2  5'b00001
`define ALU_SUB_2  5'b00010

`endif // ALU_VH
